
module ALU(



    
)